netcdf q {
dimensions:
	Layer = 45 ;
variables:
	double Layer(Layer) ;
		Layer:long_name = "Layer Target Potential Density" ;
		Layer:units = "kg m-3" ;
		Layer:cartesian_axis = "Z" ;
		Layer:positive = "up" ;

// global attributes:
		:filename = "coordinate_nk45.nc" ;

data:

   Layer = 1022.6, 1022.81, 1023.07, 1023.32, 1023.56, 1023.79, 1024.0, 1024.21, 1024.41, 1024.59, 1024.77, 1024.94, 1025.13, 1025.36, 1025.56, 1025.75, 1025.94, 1026.1, 1026.25, 1026.4, 1026.54, 1026.65, 1026.77, 1026.88, 1026.97, 1027.07, 1027.18, 1027.29, 1027.37, 1027.46, 1027.54, 1027.61, 1027.66, 1027.71, 1027.77, 1027.82, 1027.85, 1027.89, 1027.94, 1027.99, 1028.02, 1028.05, 1028.08, 1028.09, 1028.1;

}
